//////////////////////////////////////////////////////////////////////////////////
// 
// Create Date:    13:34:31 10/22/2019 
// Design Name: 	 Ferney alberto Beltran Molina
// Module Name:    VGA_Driver 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module VGA_Driver640x480 (
	input rst,
	input clk, 				// 25MHz  para 60 hz de 640x480
	input  [7:0] pixelIn, 	// entrada del valor de color  pixel 
	
	output  [7:0] pixelOut, // salida del valor pixel a la VGA 
	output  Hsync_n,		// seÃ±al de sincronizaciÃ³n en horizontal negada
	output  Vsync_n,		// seÃ±al de sincronizaciÃ³n en vertical negada 
	output  [9:0] posX, 	// posicion en horizontal del pixel siguiente
	output  [8:0] posY 		// posicion en vertical  del pixel siguiente
);

//parámetros
localparam SCREEN_X = 640; 	// tamaño de la pantalla visible en horizontal 
localparam FRONT_PORCH_X =16;  // margen superior
localparam SYNC_PULSE_X = 96;  // hsync length
localparam BACK_PORCH_X = 48;  //margen inferior
localparam TOTAL_SCREEN_X = SCREEN_X + FRONT_PORCH_X + SYNC_PULSE_X + BACK_PORCH_X; 	// total pixel pantalla en horizontal (800)


localparam SCREEN_Y = 480; 	// tamaño de la pantalla visible en Vertical 
localparam FRONT_PORCH_Y = 10;  //margen superior
localparam SYNC_PULSE_Y = 2;   //Vsync length
localparam BACK_PORCH_Y = 33;  //margen inferior
localparam TOTAL_SCREEN_Y = SCREEN_Y + FRONT_PORCH_Y + SYNC_PULSE_Y + BACK_PORCH_Y; 	// total pixel pantalla en Vertical (525)

//registros
reg  [9:0] countX;
reg  [8:0] countY;

//asignaciones (combinacional)
assign posX = countX;
assign posY = countY;

assign pixelOut = (countX < SCREEN_X) ? (pixelIn) : (8'b00000000);

assign Hsync_n = ~((countX >= SCREEN_X + FRONT_PORCH_X) && (countX < SCREEN_X + FRONT_PORCH_X + SYNC_PULSE_X)); 
assign Vsync_n = ~((countY >= SCREEN_Y + FRONT_PORCH_Y) && (countY < SCREEN_Y + FRONT_PORCH_Y + SYNC_PULSE_Y));

//logica contadores
always @(posedge clk) begin
	if (rst) begin
		countX <= 10'b0;
		countY <= 10'b0;
	end
	else begin 
		if (countX >= (TOTAL_SCREEN_X - 1)) begin
			countX <= 0;
			if (countY >= (TOTAL_SCREEN_Y - 1)) begin
				countY <= 0;
			end 
			else begin
				countY <= countY + 1;
			end
		end 
		else begin
			countX <= countX + 1;
			countY <= countY;
		end
	end
end

endmodule
